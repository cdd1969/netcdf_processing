netcdf cut_stitched {
dimensions:
	getmGrid3D_getm_1 = 139 ;
	getmGrid2D_getm_1 = 139 ;
	getmGrid2D_getm_2 = 98 ;
	getmGrid3D_getm_2 = 98 ;
	pelagic_horizontal_grid_2 = 14 ;
	pelagic_horizontal_grid_1 = 14 ;
	time = 37 ;
	getmGrid3D_getm_3 = 2 ;
variables:
	int getmGrid2D_getm_X(getmGrid2D_getm_1) ;
		getmGrid2D_getm_X:units = "1" ;
		getmGrid2D_getm_X:missing_value = -1 ;
		getmGrid2D_getm_X:axis = "X" ;
	int getmGrid2D_getm_Y(getmGrid2D_getm_2) ;
		getmGrid2D_getm_Y:units = "1" ;
		getmGrid2D_getm_Y:missing_value = -1 ;
		getmGrid2D_getm_Y:axis = "Y" ;
	double getmGrid2D_getm_lat(getmGrid2D_getm_2, getmGrid2D_getm_1) ;
		getmGrid2D_getm_lat:standard_name = "latitude" ;
		getmGrid2D_getm_lat:long_name = "getmGrid2D_getm_lat" ;
		getmGrid2D_getm_lat:units = "degrees_north" ;
		getmGrid2D_getm_lat:missing_value = -990. ;
		getmGrid2D_getm_lat:formula_terms = "" ;
		getmGrid2D_getm_lat:horizontal_stagger_location = "center" ;
		getmGrid2D_getm_lat:creator = "getm" ;
	double getmGrid2D_getm_lon(getmGrid2D_getm_2, getmGrid2D_getm_1) ;
		getmGrid2D_getm_lon:standard_name = "longitude" ;
		getmGrid2D_getm_lon:long_name = "getmGrid2D_getm_lon" ;
		getmGrid2D_getm_lon:units = "degrees_east" ;
		getmGrid2D_getm_lon:missing_value = -990. ;
		getmGrid2D_getm_lon:formula_terms = "" ;
		getmGrid2D_getm_lon:horizontal_stagger_location = "center" ;
		getmGrid2D_getm_lon:creator = "getm" ;
	int getmGrid3D_getm_X(getmGrid3D_getm_1) ;
		getmGrid3D_getm_X:units = "1" ;
		getmGrid3D_getm_X:missing_value = -1 ;
		getmGrid3D_getm_X:axis = "X" ;
	int getmGrid3D_getm_Y(getmGrid3D_getm_2) ;
		getmGrid3D_getm_Y:units = "1" ;
		getmGrid3D_getm_Y:missing_value = -1 ;
		getmGrid3D_getm_Y:axis = "Y" ;
	double getmGrid3D_getm_lat(getmGrid3D_getm_2, getmGrid3D_getm_1) ;
		getmGrid3D_getm_lat:standard_name = "latitude" ;
		getmGrid3D_getm_lat:long_name = "getmGrid3D_getm_lat" ;
		getmGrid3D_getm_lat:units = "degrees_north" ;
		getmGrid3D_getm_lat:missing_value = -990. ;
		getmGrid3D_getm_lat:formula_terms = "" ;
		getmGrid3D_getm_lat:horizontal_stagger_location = "center" ;
		getmGrid3D_getm_lat:creator = "getm" ;
	double getmGrid3D_getm_lon(getmGrid3D_getm_2, getmGrid3D_getm_1) ;
		getmGrid3D_getm_lon:standard_name = "longitude" ;
		getmGrid3D_getm_lon:long_name = "getmGrid3D_getm_lon" ;
		getmGrid3D_getm_lon:units = "degrees_east" ;
		getmGrid3D_getm_lon:missing_value = -990. ;
		getmGrid3D_getm_lon:formula_terms = "" ;
		getmGrid3D_getm_lon:horizontal_stagger_location = "center" ;
		getmGrid3D_getm_lon:creator = "getm" ;
	double pelagic_horizontal_grid_lat(pelagic_horizontal_grid_2, pelagic_horizontal_grid_1) ;
		pelagic_horizontal_grid_lat:standard_name = "latitude" ;
		pelagic_horizontal_grid_lat:long_name = "pelagic_horizontal_grid_lat" ;
		pelagic_horizontal_grid_lat:units = "degree" ;
		pelagic_horizontal_grid_lat:missing_value = -990. ;
		pelagic_horizontal_grid_lat:formula_terms = "" ;
		pelagic_horizontal_grid_lat:horizontal_stagger_location = "center" ;
	double pelagic_horizontal_grid_lon(pelagic_horizontal_grid_2, pelagic_horizontal_grid_1) ;
		pelagic_horizontal_grid_lon:standard_name = "longitude" ;
		pelagic_horizontal_grid_lon:long_name = "pelagic_horizontal_grid_lon" ;
		pelagic_horizontal_grid_lon:units = "degree" ;
		pelagic_horizontal_grid_lon:missing_value = -990. ;
		pelagic_horizontal_grid_lon:formula_terms = "" ;
		pelagic_horizontal_grid_lon:horizontal_stagger_location = "center" ;
	float shear_stress_at_soil_surface(time, getmGrid2D_getm_2, getmGrid2D_getm_1) ;
		shear_stress_at_soil_surface:_FillValue = -1.e+30f ;
		shear_stress_at_soil_surface:creator = "erosed" ;
		shear_stress_at_soil_surface:numeric_precision = "NF90_REAL" ;
		shear_stress_at_soil_surface:standard_name = "shear_stress_at_soil_surface" ;
		shear_stress_at_soil_surface:long_name = "shear_stress_at_soil_surface" ;
		shear_stress_at_soil_surface:coordinates = "getmGrid2D_getm_lat getmGrid2D_getm_lon" ;
		shear_stress_at_soil_surface:missing_value = -1.e+30f ;
	double time(time) ;
		time:units = "seconds since 2002-01-01 00:00:00" ;
		time:standard_name = "time" ;
	float water_depth_at_soil_surface(time, getmGrid2D_getm_2, getmGrid2D_getm_1) ;
		water_depth_at_soil_surface:_FillValue = -1.e+30f ;
		water_depth_at_soil_surface:units = "m" ;
		water_depth_at_soil_surface:creator = "getm" ;
		water_depth_at_soil_surface:numeric_precision = "NF90_REAL" ;
		water_depth_at_soil_surface:standard_name = "water_depth_at_soil_surface" ;
		water_depth_at_soil_surface:long_name = "water_depth_at_soil_surface" ;
		water_depth_at_soil_surface:coordinates = "getmGrid2D_getm_lat getmGrid2D_getm_lon" ;
		water_depth_at_soil_surface:missing_value = -1.e+30f ;
	float concentration_of_SPM_in_water_001(time, getmGrid3D_getm_3, getmGrid3D_getm_2, getmGrid3D_getm_1) ;
		concentration_of_SPM_in_water_001:_FillValue = -1.e+30f ;
		concentration_of_SPM_in_water_001:creator = "fabm_pelagic" ;
		concentration_of_SPM_in_water_001:units = "mg/l" ;
		concentration_of_SPM_in_water_001:mean_particle_diameter = 1.5e-05 ;
		concentration_of_SPM_in_water_001:particle_density = 1200. ;
		concentration_of_SPM_in_water_001:external_index = 3 ;
		concentration_of_SPM_in_water_001:numeric_precision = "NF90_REAL" ;
		concentration_of_SPM_in_water_001:standard_name = "concentration_of_SPM_in_water" ;
		concentration_of_SPM_in_water_001:long_name = "concentration_of_SPM_in_water" ;
		concentration_of_SPM_in_water_001:coordinates = "getmGrid3D_getm_level getmGrid3D_getm_lat getmGrid3D_getm_lon" ;
		concentration_of_SPM_in_water_001:missing_value = -1.e+30f ;
	float concentration_of_SPM_in_water_002(time, getmGrid3D_getm_3, getmGrid3D_getm_2, getmGrid3D_getm_1) ;
		concentration_of_SPM_in_water_002:_FillValue = -1.e+30f ;
		concentration_of_SPM_in_water_002:creator = "fabm_pelagic" ;
		concentration_of_SPM_in_water_002:units = "mg/l" ;
		concentration_of_SPM_in_water_002:mean_particle_diameter = 1.e-05 ;
		concentration_of_SPM_in_water_002:particle_density = 1200. ;
		concentration_of_SPM_in_water_002:external_index = 2 ;
		concentration_of_SPM_in_water_002:numeric_precision = "NF90_REAL" ;
		concentration_of_SPM_in_water_002:standard_name = "concentration_of_SPM_in_water" ;
		concentration_of_SPM_in_water_002:long_name = "concentration_of_SPM_in_water" ;
		concentration_of_SPM_in_water_002:coordinates = "getmGrid3D_getm_level getmGrid3D_getm_lat getmGrid3D_getm_lon" ;
		concentration_of_SPM_in_water_002:missing_value = -1.e+30f ;
	float concentration_of_SPM_in_water_003(time, getmGrid3D_getm_3, getmGrid3D_getm_2, getmGrid3D_getm_1) ;
		concentration_of_SPM_in_water_003:_FillValue = -1.e+30f ;
		concentration_of_SPM_in_water_003:creator = "fabm_pelagic" ;
		concentration_of_SPM_in_water_003:units = "mg/l" ;
		concentration_of_SPM_in_water_003:mean_particle_diameter = 4.e-05 ;
		concentration_of_SPM_in_water_003:particle_density = 1200. ;
		concentration_of_SPM_in_water_003:external_index = 1 ;
		concentration_of_SPM_in_water_003:numeric_precision = "NF90_REAL" ;
		concentration_of_SPM_in_water_003:standard_name = "concentration_of_SPM_in_water" ;
		concentration_of_SPM_in_water_003:long_name = "concentration_of_SPM_in_water" ;
		concentration_of_SPM_in_water_003:coordinates = "getmGrid3D_getm_level getmGrid3D_getm_lat getmGrid3D_getm_lon" ;
		concentration_of_SPM_in_water_003:missing_value = -1.e+30f ;
	double getmGrid3D_getm_layer(getmGrid3D_getm_3, getmGrid3D_getm_2, getmGrid3D_getm_1) ;
		getmGrid3D_getm_layer:standard_name = "layer" ;
		getmGrid3D_getm_layer:long_name = "getmGrid3D_getm_layer" ;
		getmGrid3D_getm_layer:units = "1" ;
		getmGrid3D_getm_layer:missing_value = -990. ;
		getmGrid3D_getm_layer:formula_terms = "" ;
		getmGrid3D_getm_layer:horizontal_stagger_location = "center" ;
		getmGrid3D_getm_layer:creator = "getm" ;
}
